--------------------------------------------------------------------------------
-- Company: Fermilab
-- Engineer: Collin Bradford
--
-- Create Date:   11:31:15 06/17/2016
-- Design Name:   
-- Module Name:   D:/cbradford/RegisterSet-2.0/GEL_CAPTAN/throttle_tb.vhd
-- Project Name:  dig_mac
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: throttle
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY throttle_tb IS
END throttle_tb;
 
ARCHITECTURE behavior OF throttle_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT throttle
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         throttle : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '1';

 	--Outputs
   signal throttley : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: throttle PORT MAP (
          clk => clk,
          rst => rst,
          throttle => throttley
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		rst <= '0';

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
