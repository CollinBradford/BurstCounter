--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:06:57 06/01/2016
-- Design Name:   
-- Module Name:   D:/cbradford/MainProjectRegisterSet/GEL_CAPTAN/WriteRegister_tb.vhd
-- Project Name:  dig_mac
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: WriteRegistser
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY WriteRegister_tb IS
END WriteRegister_tb;
 
ARCHITECTURE behavior OF WriteRegister_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT WriteRegistser
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         rx_addr : IN  std_logic_vector(31 downto 0);
         rx_data : IN  std_logic_vector(63 downto 0);
         rx_wren : IN  std_logic;
         user_ready : OUT  std_logic;
         reg_out : OUT  std_logic_vector(63 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '1';
   signal clk : std_logic := '0';
   signal rx_addr : std_logic_vector(31 downto 0) := (others => '0');
   signal rx_data : std_logic_vector(63 downto 0) := (others => '0');
   signal rx_wren : std_logic := '0';

 	--Outputs
   signal user_ready : std_logic;
   signal reg_out : std_logic_vector(63 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: WriteRegistser PORT MAP (
          rst => rst,
          clk => clk,
          rx_addr => rx_addr,
          rx_data => rx_data,
          rx_wren => rx_wren,
          user_ready => user_ready,
          reg_out => reg_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		rst <= '0';

      wait for clk_period * 9;
		
		rx_data <= (others => '1');
		rx_wren <= '1';
		
		wait for clk_period * 3;
		
		rx_data <= (others => '0');
		rx_wren <= '0';

      wait;
   end process;

END;
